`timescale 1s/100ms
`include "comparator4.v"

module comparator4_tb();
	reg [0:3]a;
	reg [0:3]b;
	wire g;
	wire e;
	wire l;

	comparator4 myComparator(a, b, g, e, l);

	initial
	begin 
		$monitor("a = %4b, b = %4b, g = %b, e = %b, l = %b", a, b, g, e, l);
		$dumpfile ("comparator4.vcd");
		$dumpvars (0, comparator4_tb);
		a = 4'b0000; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b0001; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b0010; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b0011; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b0100; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b0101; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b0110; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b0111; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b1000; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b1001; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b1010; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b1011; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b1100; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b1101; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b1110; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;

		a = 4'b1111; b = 4'b0000; #1;
		b = 4'b0001; #1;
		b = 4'b0010; #1;
		b = 4'b0011; #1;
		b = 4'b0100; #1;
		b = 4'b0101; #1;
		b = 4'b0110; #1;
		b = 4'b0111; #1;
		b = 4'b1000; #1;
		b = 4'b1001; #1;
		b = 4'b1010; #1;
		b = 4'b1011; #1;
		b = 4'b1100; #1;
		b = 4'b1101; #1;
		b = 4'b1110; #1;
		b = 4'b1111; #1;
		$finish;
	end
endmodule